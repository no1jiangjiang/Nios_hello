// hello.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module hello (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
